LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--端口定义
ENTITY LED_DISP IS
	PORT(
		IND:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		LEDN:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		
		SEG:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTD:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY LED_DISP;

--实体描述
ARCHITECTURE ART OF LED_DISP IS

SIGNAL IND:STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL  

SIGNAL s_SEG: STD_LOGIC_VECTOR(7 DOWNTO 0) ;
SIGNAL s_OUTD: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
P1: PROCESS(CLK,RST) IS
BEGIN
	IF(CLK'EVENT AND CLK='1') THEN
	END IF;
END PROCESS P1;
P2:	PROCESS(LEDN,IND) IS
	BEGIN
		CASE LEDN IS
			WHEN "000"=>s_SEG<="00000001";
			WHEN "001"=>s_SEG<="00000010";
			WHEN "010"=>s_SEG<="00000100";
			WHEN "011"=>s_SEG<="00001000";
			WHEN "100"=>s_SEG<="00010000";
			WHEN "101"=>s_SEG<="00100000";
			WHEN "110"=>s_SEG<="01000000";
			WHEN "111"=>s_SEG<="10000000";
			WHEN OTHERS =>s_SEG<="XXXXXXXX";
		END CASE;
		CASE IND IS
			WHEN "0000" => s_OUTD <= "11000000";
			WHEN "0001" => s_OUTD <= "11111001"; 
			WHEN "0010" => s_OUTD <= "10100100"; 
			WHEN "0011" => s_OUTD <= "10110000";
			
			WHEN "0100" => s_OUTD <= "10011001"; 
			WHEN "0101" => s_OUTD <= "10010010"; 
			WHEN "0110" => s_OUTD <= "10000010"; 
			WHEN "0111" => s_OUTD <= "11111000";
			
			WHEN "1000" => s_OUTD <= "10000000";
			WHEN "1001" => s_OUTD <= "10010000"; 
			WHEN "1010" => s_OUTD <= "10001000"; 
			WHEN "1011" => s_OUTD <= "10000011";
			
			WHEN "1100" => s_OUTD <= "11000110"; 
			WHEN "1101" => s_OUTD <= "10100001"; 
			WHEN "1110" => s_OUTD <= "10000110"; 
			WHEN "1111" => s_OUTD <= "10001110";
			WHEN OTHERS => s_OUTD <= "XXXXXXXX";
		END CASE;		
	END PROCESS P2;
	
SEG<=s_SEG;
OUTD<=s_OUTD;	
END ARCHITECTURE ART;
	