LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TOP IS
	PORT(
	I:STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY TOP;

ARCHITECTURE ART OF TOP IS
BEGIN

END ARCHITECTURE ART;

	