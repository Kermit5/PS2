LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--实体定义
ENTITY DATA_SCAN IS
	PORT(
		SYS_CLK,K_DATA,K_CLOCK,RST:IN STD_LOGIC;
		DATA:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		PA:INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		ZHJS:INOUT STD_LOGIC
	);
END ENTITY DATA_SCAN;

ARCHITECTURE ART OF DATA_SCAN IS
--信号定义
SIGNAL TEMP:STD_LOGIC_VECTOR(11 DOWNTO 0):="000000000000";

SIGNAL CUR_KBCLK,PRE_KBCLK:STD_LOGIC;
--开始信号
SIGNAL START:STD_LOGIC;
--使能信号
SIGNAL EN:STD_LOGIC;
--计数变量
SIGNAL CNT:STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN

P1: PROCESS(SYS_CLK,RST) IS
	BEGIN
		IF(RST='0') THEN
			ZHJS<='0';
			CNT<="0000";
			START<='0';
		ELSE
			IF(SYS_CLK'EVENT AND SYS_CLK='1') THEN
				PRE_KBCLK<=CUR_KBCLK;
				CUR_KBCLK<=K_CLOCK;
				--采样数据，一共12位，1位起始位，8位数据位，1位校验位，1位结束位
				IF(PRE_KBCLK>CUR_KBCLK) THEN
					CASE CNT IS 
						WHEN "0000" => TEMP(0)<=K_DATA;
						WHEN "0001" => TEMP(1)<=K_DATA;
						WHEN "0010" => TEMP(2)<=K_DATA;
						WHEN "0011" => TEMP(3)<=K_DATA;
						
						WHEN "0100" => TEMP(4)<=K_DATA;
						WHEN "0101" => TEMP(5)<=K_DATA;
						WHEN "0110" => TEMP(6)<=K_DATA;
						WHEN "0111" => TEMP(7)<=K_DATA;
						
						WHEN "1000" => TEMP(8)<=K_DATA;
						WHEN "1001" => TEMP(9)<=K_DATA;
						WHEN "1010" => TEMP(10)<=K_DATA;
						WHEN "1011" => TEMP(11)<=K_DATA;
						
						WHEN OTHERS => TEMP(0)<='X';
					END CASE;
					--数据接收完成
					IF(CNT="1010") THEN
						ZHJS<='0';
					ELSE
						ZHJS<='1';
					END IF;
					IF(CNT="1011") THEN
						CNT<="0001";
					ELSE
						CNT<=CNT+'1';
					END IF; 	
				END IF;
				IF(CNT>"0001" AND CNT<"1010") THEN
					START<='1';
				ELSE
					START<='0';
				END IF;
			END IF;
		END IF;
END PROCESS P1;


P2: PROCESS(SYS_CLK) IS
BEGIN
	IF(SYS_CLK'EVENT AND SYS_CLK='1') THEN
		IF(START='1') THEN
			PA<="00000000";
		ELSE
			PA<=TEMP(9 DOWNTO 2);
		END IF;
		IF(ZHJS='0') THEN
			DATA<=PA;
		END IF;
	END IF;
END PROCESS P2;
END ARCHITECTURE ART;

